* Generator created 01 Oct 2022 by John Lutz. Editeded 02 Oct 2022
* This file generated on: 02 Oct 2022

.SUBCKT ring_osc_1 in0 out12 vdd 0

    x0 in0 out0 vdd 0 inverter params:
    + tplv=0.0721u tpotv=2.0344n tpwv=236.1375n 
    + tnln=0.072u tnwn=134.4984n tnotv=1.7233n 

    x1 out0 out1 vdd 0 inverter params:
    + tplv=0.0655u tpotv=2.1131n tpwv=194.5286n 
    + tnln=0.0618u tnwn=133.4563n tnotv=1.95n 

    x2 out1 out2 vdd 0 inverter params:
    + tplv=0.0675u tpotv=1.7714n tpwv=249.9654n 
    + tnln=0.0679u tnwn=128.8598n tnotv=1.7361n 

    x3 out2 out3 vdd 0 inverter params:
    + tplv=0.0679u tpotv=1.8464n tpwv=231.259n 
    + tnln=0.0737u tnwn=134.0122n tnotv=1.8945n 

    x4 out3 out4 vdd 0 inverter params:
    + tplv=0.0592u tpotv=1.7675n tpwv=204.9133n 
    + tnln=0.0625u tnwn=136.4309n tnotv=1.7493n 

    x5 out4 out5 vdd 0 inverter params:
    + tplv=0.0745u tpotv=1.772n tpwv=201.9264n 
    + tnln=0.0684u tnwn=136.6653n tnotv=1.7413n 

    x6 out5 out6 vdd 0 inverter params:
    + tplv=0.0659u tpotv=2.0613n tpwv=232.2619n 
    + tnln=0.0735u tnwn=126.6155n tnotv=1.7719n 

    x7 out6 out7 vdd 0 inverter params:
    + tplv=0.0739u tpotv=2.0528n tpwv=204.2462n 
    + tnln=0.0612u tnwn=130.6029n tnotv=1.9697n 

    x8 out7 out8 vdd 0 inverter params:
    + tplv=0.0743u tpotv=2.1433n tpwv=199.8904n 
    + tnln=0.0735u tnwn=137.3065n tnotv=2.0074n 

    x9 out8 out9 vdd 0 inverter params:
    + tplv=0.0616u tpotv=1.9421n tpwv=226.7772n 
    + tnln=0.0715u tnwn=121.0625n tnotv=1.7217n 

    x10 out9 out10 vdd 0 inverter params:
    + tplv=0.0696u tpotv=1.7732n tpwv=224.1744n 
    + tnln=0.0569u tnwn=129.0007n tnotv=1.7176n 

    x11 out10 out11 vdd 0 inverter params:
    + tplv=0.0704u tpotv=1.9575n tpwv=250.3129n 
    + tnln=0.0712u tnwn=135.4386n tnotv=1.9944n 

    x12 out11 out12 vdd 0 inverter params:
    + tplv=0.0701u tpotv=2.0098n tpwv=231.0229n 
    + tnln=0.0601u tnwn=113.7579n tnotv=1.9029n 

.ENDS ring_osc.end
