* Generator created 01 Oct 2022 by John Lutz. Editeded 02 Oct 2022
* This file generated on: 02 Oct 2022

.SUBCKT ring_osc_5 in0 out12 vdd 0

    x0 in0 out0 vdd 0 inverter params:
    + tplv=0.0646u tpotv=1.9972n tpwv=232.3163n 
    + tnln=0.0655u tnwn=149.1682n tnotv=1.9773n 

    x1 out0 out1 vdd 0 inverter params:
    + tplv=0.0669u tpotv=2.0127n tpwv=205.5075n 
    + tnln=0.064u tnwn=117.1927n tnotv=1.8932n 

    x2 out1 out2 vdd 0 inverter params:
    + tplv=0.0701u tpotv=2.0878n tpwv=219.2931n 
    + tnln=0.0737u tnwn=138.2593n tnotv=1.8959n 

    x3 out2 out3 vdd 0 inverter params:
    + tplv=0.0708u tpotv=2.0442n tpwv=194.5407n 
    + tnln=0.07u tnwn=113.343n tnotv=1.9532n 

    x4 out3 out4 vdd 0 inverter params:
    + tplv=0.0683u tpotv=1.8968n tpwv=238.8489n 
    + tnln=0.0577u tnwn=148.4908n tnotv=1.7123n 

    x5 out4 out5 vdd 0 inverter params:
    + tplv=0.0634u tpotv=1.9893n tpwv=219.927n 
    + tnln=0.0736u tnwn=141.1634n tnotv=1.8454n 

    x6 out5 out6 vdd 0 inverter params:
    + tplv=0.0731u tpotv=2.0539n tpwv=201.1739n 
    + tnln=0.0715u tnwn=120.6058n tnotv=1.844n 

    x7 out6 out7 vdd 0 inverter params:
    + tplv=0.0657u tpotv=2.0434n tpwv=233.9119n 
    + tnln=0.0705u tnwn=122.541n tnotv=1.8113n 

    x8 out7 out8 vdd 0 inverter params:
    + tplv=0.0747u tpotv=1.788n tpwv=202.8024n 
    + tnln=0.0705u tnwn=147.0969n tnotv=1.9816n 

    x9 out8 out9 vdd 0 inverter params:
    + tplv=0.0712u tpotv=2.1286n tpwv=235.028n 
    + tnln=0.0698u tnwn=144.1824n tnotv=1.9458n 

    x10 out9 out10 vdd 0 inverter params:
    + tplv=0.0732u tpotv=1.8502n tpwv=186.9993n 
    + tnln=0.071u tnwn=137.3481n tnotv=1.8065n 

    x11 out10 out11 vdd 0 inverter params:
    + tplv=0.0698u tpotv=1.9654n tpwv=209.3332n 
    + tnln=0.0604u tnwn=130.6278n tnotv=1.8869n 

    x12 out11 out12 vdd 0 inverter params:
    + tplv=0.0594u tpotv=1.8337n tpwv=231.8177n 
    + tnln=0.0563u tnwn=119.0337n tnotv=1.7495n 

.ENDS ring_osc.end
